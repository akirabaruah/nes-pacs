module nes ();

endmodule
